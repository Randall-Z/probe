 RL CIRCUIT AND PROBE
 VS 1 0 SIN(0 10 100 0 0 0 )
 L1 1 2 1MH
 R1 2 1 100
 *CONTROL STATEMENT
 .TRAN 1.0E-3 3.0E-2
 .PROBE.END